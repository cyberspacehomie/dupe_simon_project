// Nothing goes in this module
// just module instances and the state machine!
module top(
	


);

endmodule
