// Nothing goes in this module
// just module instances!
module top(
	);

endmodule
